module test();
import pkg::*;
  porsche p_h;
  initial begin
    p_h = new();
  end
endmodule: test